*-----------------------------------------------------------------------------
*
* To use a subcircuit, the name must begin with 'X'.  For example:
* X1 1 2 3 4 5 uA741
*
* connections:   non-inverting input
*                |  inverting input
*                |  |  positive power supply
*                |  |  |  negative power supply
*                |  |  |  |  output
*                |  |  |  |  |
.subckt uA741    1  2  3  4  5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends



.options savecurrents

Vcc vcc 0 5.0
Vee vee 0 -5.0
Vin in 0 0

X1 inv_out inv_in vcc vee outb uA741


*R1 and C1
C1 in inv_in 220n
R1 inv_in 0 1k


*R2 and C2
R2 outb out 1k
C2 out 0 110n

*R3 and R4 fixed
R3 inv_out outb 120k
R4 inv_out 0 1k


Vout out 0 0 ac 1 sin(0 1 1000)

.op
.end

.control

print all

* frequency analysis
ac dec 10 10 100MEG

*MEASURE
*output impedance in kohm
let outputimpedance = -(v(out)[20]/Vout#branch[20])

echo "outimpedance_TAB"
print outputimpedance
echo "outimpedance_END"


.endc 

