*
* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents

*Circuit description

.INCLUDE sim2data.cir

*.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "****************"
echo  "Operating point"
echo "****************"

echo  "op2_TAB"
print all
echo  "op2_END"

quit
.endc

.end
