*
* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents

*Voltage source

Vs n1 0 0
V0 n7 n9 DC 0

*Voltage source in the place of Capacitor (v6-v8)

Vx n8 n6 8.49302

*Dependent Sources

H0 n5 n8 V0 8.36641247715k
G0 n6 n3 n2 n5 7.28209304852m

* Resistors

R1 n1 n2 1.04765357286k
R2 n3 n2 2.06140068334k
R3 n2 n5 3.03459085363k
R4 n5 0 4.00398818216k
R5 n5 n6 3.11499853456k 
R6 0 n7 2.04588646991k
R7 n9 n8 1.04390152967k

*.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "****************"
echo  "Operating point"
echo "****************"

echo  "op_TAB"
print all
echo  "op_END"

quit
.endc

.end
