*
* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents

*Circuit description

*AC In and transformer description
VIN n1 0 SIN(0 230 50 0 0)
F1 n1 0 E2 17
E2 n2 0 n1 0 0.058824

*Envelope Detector
R1 n2 n3 50k
C1 n3 0 1u
D1 n3 n4 Default
D2 n4 n5 Default
D3 n5 0 Default
D6 0 n6 Default
D7 n6 n7 Default
D8 n7 n3 Default
R2 n3 0 1k
C2 n3 0 1u 

*Voltage Regulator


.model Default D
*.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "****************"
echo  "Operating point"
echo "****************"

echo  "op1_TAB"
print all
echo  "op1_END"

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 2e-1

hardcopy transientalt.ps v(n3)
echo transientalt_FIG

quit
.endc

.end
