*
* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents

*Circuit description

*AC In and transformer description
VIN n1 0 SIN(0 230 50 0 0)
F1 n1 0 E2 14
E2 n2 0 n1 0 0.071429

*Diodos manhosos
D5 n2 n7 Default
D6 0 n7 Default
D7 n8 0 Default
D8 n8 2 Default

*Envelope Detector
R1 n7 n8 50k
C0 n7 n8 10u

*Voltage Regulator
R2 n7 n4 5k
D2 n4 n5 Default
D3 n5 n6 Default
D4 n6 n9 Default
D9 n9 n10 Default
D10 n10 n11 Default
D11 n11 n12 Default
D12 n12 n13 Default
D13 n13 n14 Default
D14 n14 n15 Default
D15 n15 n16 Default
D16 n16 n17 Default
D17 n17 n18 Default
D18 n18 n19 Default
D19 n19 n20 Default
D20 n20 n21 Default
D21 n21 n22 Default
D22 n22 n23 Default
D23 n23 n24 Default
D24 n24 n8 Default
*D25 n25 n8 Default

*Calculate Values
*ripple = max(v(n4)-v(n8)) - min(v(n4)-v(n8))
*average = avg(v(n4)-v(n8))

.model Default D
*.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "****************"
echo  "Operating point"
echo "****************"

echo  "op1_TAB"
print all
echo  "op1_END"

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 5e-5 2e-1

hardcopy transientfinal.ps v(n4)-v(n8)
echo transientfinal_FIG

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 5e-5 2e-1

hardcopy transientenvelope.ps v(n7)-v(n8)
echo transientenvelope_FIG

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 5e-5 2e-1

hardcopy transient5.ps v(n4)-v(n8)-12
echo transient5_FIG

quit
.endc

.end
