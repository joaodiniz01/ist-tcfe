*
* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents

*Circuit description

.INCLUDE sim3data.cir

*.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

*echo "****************"
*echo  "Operating point"
*echo "****************"

*echo  "op_TAB"
*print all
*echo  "op_END"

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-3 20e-3

hardcopy ../doc/transient3.ps v(n6)
echo transient3_FIG


quit
.endc

.end
